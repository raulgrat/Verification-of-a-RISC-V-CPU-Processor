/* DISCLAIMER:

This file is intentionally left blank here for whichever testbench you would like to run.
Simply just paste the corresponding Testbench file into this testbench.sv and change the first line of the files.f to corresponding design.
Alternatively, this page can be left blank and to run the specific testbench, you may change the second line of the files.f to the corresponding testbench file

***Be sure to check Use run.bash shell script***

The testbenches we made were used for verifying the individual module components of the RISCV CPU


This verification project was done by the following members:
- Jack Gao
- Francisco Soriano
- Raul Graterol Medina

*/
